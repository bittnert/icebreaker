module uart_rx (input CLK, input rst, output rx_ready, output[7:0] rx_data);


endmodule

